module axi_cov_top;
  //Define the interface hierarchy
  `define axi_if dut_top
  //Checker connection
  axi_cov axi_cov();
    // defparam axi_cov.INST_NAME = "AXI_FUNCTIONAL_COVERAGE";
    assign axi_cov.aclk    = `axi_if.aclk;
    assign axi_cov.aresetn = `axi_if.aresetn;
    assign axi_cov.awvalid = `axi_if.awvalid;
    assign axi_cov.awready = `axi_if.awready;
    assign axi_cov.awid    = `axi_if.awid;
    assign axi_cov.awaddr  = `axi_if.awaddr;
    assign axi_cov.awlen   = `axi_if.awlen;
    assign axi_cov.awsize  = `axi_if.awsize;
    assign axi_cov.awburst = `axi_if.awburst;
    assign axi_cov.wvalid  = `axi_if.wvalid;
    assign axi_cov.wdata   = `axi_if.wdata;
    assign axi_cov.wstrb   = `axi_if.wstrb;
    assign axi_cov.wlast   = `axi_if.wlast;
    assign axi_cov.wready  = `axi_if.wready;
    assign axi_cov.bready  = `axi_if.bready;
    assign axi_cov.bvalid  = `axi_if.bvalid;
    assign axi_cov.bresp  = `axi_if.bresp;
    assign axi_cov.bid  = `axi_if.bid;
    assign axi_cov.arvalid = `axi_if.arvalid;
    assign axi_cov.arready = `axi_if.arready;
    assign axi_cov.arid    = `axi_if.arid;
    assign axi_cov.araddr  = `axi_if.araddr;
    assign axi_cov.arlen   = `axi_if.arlen;
    assign axi_cov.arsize  = `axi_if.arsize;
    assign axi_cov.arburst = `axi_if.arburst;
    assign axi_cov.rvalid  = `axi_if.rvalid;
    assign axi_cov.rdata   = `axi_if.rdata;
    assign axi_cov.rlast   = `axi_if.rlast;
    assign axi_cov.rready  = `axi_if.rready;
    assign axi_cov.rresp  = `axi_if.rresp;
    assign axi_cov.rid  = `axi_if.rid;
endmodule
 